module sum3bits ();

endmodule