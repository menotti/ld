module vector(
  input [3:0] a,
  input [3:0] b,
  output [3:0] a_bitwise_or_b,
  output a_logical_or_b,
  output a_reduction_or,
  output b_reduction_or,
  output [7:0] not_a_not_b);
  // Implemente as operações para cada uma das saídas usando o modelo
  // assign a_bitwise_or_b = ... ;

endmodule
