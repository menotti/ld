module top(
	output GPIO_0_D0);	
	
	assign GPIO_0_D0 = 1'b1; 
endmodule
