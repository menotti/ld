
module top (
    input  [31:0] a,
    input  [31:0] b,
    input         sub,         // 0 = soma, 1 = subtração
    output [31:0] result,
    output        carry_out,
    output        overflow);



endmodule