module top(
  input [1:0] SW,
  output [6:0] HEX0);
  // instancie e conecte os módulos a seguir


endmodule
