module moore (
    input clk, rst, w, 
    output z);



endmodule