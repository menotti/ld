module tb_hello;
    hello dut();
endmodule 
