module top(
  input CLOCK_50,
  input [3:0] SW,
  input [1:0] KEY,
  output [3:0] f); 	//simulacao  
  //output [6:0] HEX0);	//implementacao  
  
  wire [3:0] a, b;
 


endmodule