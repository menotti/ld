module mealy (
    input clk, rst, w, 
    output z);



endmodule