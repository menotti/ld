module top (
    input a, b, c, d,
    output f1, f2, f3);



endmodule