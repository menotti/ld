module addsum4bits (
  input op,
  input signed [3:0] x, y,
  output signed [3:0] s,
  output ov);
  
  // 1. Implemente aqui o somador/subtrator aqui e simule para testar 


endmodule