// Use este modulo quando for gravar na placa
/* 
module top(
  input op, // Usar o pb[0]
  input [2:0] sw, // x
  input [2:0] ja, // y
  output [3:0] jb, // segmentos [a-d]
  output [3:0] jc); // segmentos [e-f]+cat

endmodule
*/


module addsum4bits (
  input op,
  input [3:0] x, y,
  output [3:0] s,
  output ov);
  // Implemente aqui o somador/subtrator
  
  
endmodule
