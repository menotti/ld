module hello;
    // uncomment the following lines
    //initial
    //  $display("Hello, Verilog!");
endmodule
