module top (
    input [31:0] in, 
    input [1:0] sel, 
    output [7:0] out);

    //declare os fios intermediarios 

    // instancie os muxes que precisar 



endmodule